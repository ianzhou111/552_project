module seven_decode(
    input [6:0] in,
    output reg [127:0] out
);

always @(*) begin
    case (in)
        7'h00: out = 128'h1;
        7'h01: out = 128'h2;
        7'h02: out = 128'h4;
        7'h03: out = 128'h8;
        7'h04: out = 128'h10;
        7'h05: out = 128'h20;
        7'h06: out = 128'h40;
        7'h07: out = 128'h80;
        7'h08: out = 128'h100;
        7'h09: out = 128'h200;
        7'h0A: out = 128'h400;
        7'h0B: out = 128'h800;
        7'h0C: out = 128'h1000;
        7'h0D: out = 128'h2000;
        7'h0E: out = 128'h4000;
        7'h0F: out = 128'h8000;
        7'h10: out = 128'h10000;
        7'h11: out = 128'h20000;
        7'h12: out = 128'h40000;
        7'h13: out = 128'h80000;
        7'h14: out = 128'h100000;
        7'h15: out = 128'h200000;
        7'h16: out = 128'h400000;
        7'h17: out = 128'h800000;
        7'h18: out = 128'h1000000;
        7'h19: out = 128'h2000000;
        7'h1A: out = 128'h4000000;
        7'h1B: out = 128'h8000000;
        7'h1C: out = 128'h10000000;
        7'h1D: out = 128'h20000000;
        7'h1E: out = 128'h40000000;
        7'h1F: out = 128'h80000000;
        7'h20: out = 128'h100000000;
        7'h21: out = 128'h200000000;
        7'h22: out = 128'h400000000;
        7'h23: out = 128'h800000000;
        7'h24: out = 128'h1000000000;
        7'h25: out = 128'h2000000000;
        7'h26: out = 128'h4000000000;
        7'h27: out = 128'h8000000000;
        7'h28: out = 128'h10000000000;
        7'h29: out = 128'h20000000000;
        7'h2A: out = 128'h40000000000;
        7'h2B: out = 128'h80000000000;
        7'h2C: out = 128'h100000000000;
        7'h2D: out = 128'h200000000000;
        7'h2E: out = 128'h400000000000;
        7'h2F: out = 128'h800000000000;
        7'h30: out = 128'h1000000000000;
        7'h31: out = 128'h2000000000000;
        7'h32: out = 128'h4000000000000;
        7'h33: out = 128'h8000000000000;
        7'h34: out = 128'h10000000000000;
        7'h35: out = 128'h20000000000000;
        7'h36: out = 128'h40000000000000;
        7'h37: out = 128'h80000000000000;
        7'h38: out = 128'h100000000000000;
        7'h39: out = 128'h200000000000000;
        7'h3A: out = 128'h400000000000000;
        7'h3B: out = 128'h800000000000000;
        7'h3C: out = 128'h1000000000000000;
        7'h3D: out = 128'h2000000000000000;
        7'h3E: out = 128'h4000000000000000;
        7'h3F: out = 128'h8000000000000000;
        7'h40: out = 128'h10000000000000000;
        7'h41: out = 128'h20000000000000000;
        7'h42: out = 128'h40000000000000000;
        7'h43: out = 128'h80000000000000000;
        7'h44: out = 128'h100000000000000000;
        7'h45: out = 128'h200000000000000000;
        7'h46: out = 128'h400000000000000000;
        7'h47: out = 128'h800000000000000000;
        7'h48: out = 128'h1000000000000000000;
        7'h49: out = 128'h2000000000000000000;
        7'h4A: out = 128'h4000000000000000000;
        7'h4B: out = 128'h8000000000000000000;
        7'h4C: out = 128'h10000000000000000000;
        7'h4D: out = 128'h20000000000000000000;
        7'h4E: out = 128'h40000000000000000000;
        7'h4F: out = 128'h80000000000000000000;
        7'h50: out = 128'h100000000000000000000;
        7'h51: out = 128'h200000000000000000000;
        7'h52: out = 128'h400000000000000000000;
        7'h53: out = 128'h800000000000000000000;
        7'h54: out = 128'h1000000000000000000000;
        7'h55: out = 128'h2000000000000000000000;
        7'h56: out = 128'h4000000000000000000000;
        7'h57: out = 128'h8000000000000000000000;
        7'h58: out = 128'h10000000000000000000000;
        7'h59: out = 128'h20000000000000000000000;
        7'h5A: out = 128'h40000000000000000000000;
        7'h5B: out = 128'h80000000000000000000000;
        7'h5C: out = 128'h100000000000000000000000;
        7'h5D: out = 128'h200000000000000000000000;
        7'h5E: out = 128'h400000000000000000000000;
        7'h5F: out = 128'h800000000000000000000000;
        7'h60: out = 128'h1000000000000000000000000;
        7'h61: out = 128'h2000000000000000000000000;
        7'h62: out = 128'h4000000000000000000000000;
        7'h63: out = 128'h8000000000000000000000000;
        7'h64: out = 128'h10000000000000000000000000;
        7'h65: out = 128'h20000000000000000000000000;
        7'h66: out = 128'h40000000000000000000000000;
        7'h67: out = 128'h80000000000000000000000000;
        7'h68: out = 128'h100000000000000000000000000;
        7'h69: out = 128'h200000000000000000000000000;
        7'h6a: out = 128'h400000000000000000000000000;
        7'h6b: out = 128'h800000000000000000000000000;
        7'h6c: out = 128'h1000000000000000000000000000;
        7'h6d: out = 128'h2000000000000000000000000000;
        7'h6e: out = 128'h4000000000000000000000000000;
        7'h6f: out = 128'h8000000000000000000000000000;
        7'h70: out = 128'h10000000000000000000000000000;
        7'h71: out = 128'h20000000000000000000000000000;
        7'h72: out = 128'h40000000000000000000000000000;
        7'h73: out = 128'h80000000000000000000000000000;
        7'h74: out = 128'h100000000000000000000000000000;
        7'h75: out = 128'h200000000000000000000000000000;
        7'h76: out = 128'h400000000000000000000000000000;
        7'h77: out = 128'h800000000000000000000000000000;
        7'h78: out = 128'h1000000000000000000000000000000;
        7'h79: out = 128'h2000000000000000000000000000000;
        7'h7a: out = 128'h4000000000000000000000000000000;
        7'h7b: out = 128'h8000000000000000000000000000000;
        7'h7c: out = 128'h10000000000000000000000000000000;
        7'h7d: out = 128'h20000000000000000000000000000000;
        7'h7e: out = 128'h40000000000000000000000000000000;
        7'h7f: out = 128'h80000000000000000000000000000000;
        default: out = 128'h0; 
    endcase 
end

endmodule 