module forward (output wire FwdOp1MX, output wire FwdOp1XX, output wire FwdOp2MX, output wire FwdOp2XX, input [3:0] ID_EX_Rs, input [3:0] ID_EX_Rt, input [3:0] EX_MEM_Rd, input [3:0] MEM_WB_Rd);



endmodule